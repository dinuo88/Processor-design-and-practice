/******************************************************************************
* Function: 下一程序计数器（NPC）模块
*
* 模块功能描述:
* - 此模块表示一个简单的下一程序计数器。
* - 它通过将输入的程序计数器值（pc）增加 4 个字节的偏移量来计算下一程序计数器值（npc）。
*
* 设计方法:
* - 输入的程序计数器值（pc）加上 4 用于计算下一程序计数器值（npc）。
*
******************************************************************************/

`timescale 1ns / 1ps

module NPC(
    input [31:0] pc,    // 输入的程序计数器值
    output [31:0] npc   // 输出的下一程序计数器值
);

    assign npc = pc + 32'd4;  // 下一程序计数器值等于输入值加上 4

endmodule
