/******************************************************************************
* Function: 字符串连接器（Strcat）模块
*
* 模块功能描述:
* - 此模块表示一个字符串连接器。
* - 它将一个 28 位的地址（addr28）和一个 4 位的高位（npc_high4）连接成一个 32 位的跳转地址（jump2addr）。
*
* 设计方法:
* - 使用 assign 语句将输入的高位（npc_high4）连接到输出的跳转地址（jump2addr）的高位。
* - 使用 assign 语句将输入的地址（addr28）连接到输出的跳转地址（jump2addr）的低位。
*
******************************************************************************/

`timescale 1ns / 1ps

module Strcat(
    input [27:0] addr28,        // 输入的 28 位地址
    input [3:0] npc_high4,     // 输入的 4 位高位
    
    output [31:0] jump2addr    // 输出的 32 位跳转地址
);

    assign jump2addr[31:28] = npc_high4;   // 连接输入的高位到输出的高位
    assign jump2addr[27:0] = addr28;        // 连接输入的地址到输出的低位

endmodule
