/******************************************************************************
* Function: 16位符号扩展模块
*
* 模块功能描述:
* - 此模块表示一个16位符号扩展模块，根据符号位来扩展输入为32位输出。
*
* 参数:
* - DEPTH: 输入宽度，默认为16位。
*
* 设计方法:
* - 使用一个 always 块，根据输入信号a和符号扩展信号sign_ext来进行符号扩展。
* - 如果符号扩展信号为1且输入a的符号位为1，将输出b的高16位设置为全1，其余位保持不变。
* - 否则，将输出b的高16位设置为全0，其余位保持不变。
*
******************************************************************************/

`timescale 1ns/1ps

module S_EXT16 #(parameter DEPTH = 16) (
    input [DEPTH - 1 : 0] a,     // 输入a
    input sign_ext,              // 符号扩展信号
    output reg [31 : 0] b       // 输出b
);

    always @ (a or sign_ext) begin
        if (sign_ext == 1 && a[DEPTH - 1] == 1) begin
            b[31:0] = 32'hffffffff;    // 符号扩展为全1
            b[DEPTH - 1:0] = a[DEPTH - 1:0];
        end
        else begin
            b[31:0] = 32'h00000000;    // 符号扩展为全0
            b[DEPTH - 1:0] = a[DEPTH - 1:0];
        end
    end
endmodule
